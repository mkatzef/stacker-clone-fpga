
module pll (
	clk_in_clk,
	clk_rst_reset,
	clk_out_clk);	

	input		clk_in_clk;
	input		clk_rst_reset;
	output		clk_out_clk;
endmodule
